`ifndef __MAT_MEM_TYPE__
`define __MAT_MEM_TYPE__

typedef enum {
    MAT_DATA_MEM_WRITE_DISABLE,
    MAT_DATA_MEM_WRITE_SINGLE,
    MAT_DATA_MEM_WRITE_ALL
} MatDataMemWriteOp_t;

`endif
