`default_nettype none

module MatControl
    (input logic clock,
     input logic instruction);

endmodule: MatControl
